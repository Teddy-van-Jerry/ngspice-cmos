* =============================================================================
* Circuit    : CMOS AND8 Gate Type C
* Description: AND4B * 2 + AND2 * 1
*
* Author     : Wuqiong Zhao (me@wqzhao.org)
* Date       : 2023-06-02
* License    : MIT
* =============================================================================

.title CMOS AND8C

* Parameters and Model
* -----------------------------------------------------------------------------
.param VDD='1.0V'
.temp  25
.inc ./FreePDK45/ff.inc

* Supply Voltage Source
* -----------------------------------------------------------------------------
Vdd vdd gnd VDD

* AND8B
* -----------------------------------------------------------------------------
XAND8 gnd in1 in2 in3 in4 in5 in6 in7 in8 out vdd AND8C
.inc ./and8c.inc

* Test Circuit
* -----------------------------------------------------------------------------
XTest gnd
+     ii1 ii2 ii3 ii4 ii5 ii6 ii7 ii8
+     in1 in2 in3 in4 in5 in6 in7 in8
+     out vdd               INV2_TEST
.inc ./and8_test_inv2.inc

* Input Signals
* -----------------------------------------------------------------------------
Vii1 ii1 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   3.0ns VDD
+ )

Vii2 ii2 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   3.0ns VDD
+ )

Vii3 ii3 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   3.0ns VDD
+ )

Vii4 ii4 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   3.0ns VDD
+ )

Vii5 ii5 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   3.0ns VDD
+ )

Vii6 ii6 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   3.0ns VDD
+ )

Vii7 ii7 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   3.0ns VDD
+ )

Vii8 ii8 gnd PWL
+ (
+   0.0ns  0V
+   0.9ns  0V
+   1.1ns VDD
+   1.9ns VDD
+   2.1ns  0V
+   3.0ns  0V
+ )

* Analysis
* -----------------------------------------------------------------------------
.ic    V(out)=0
.tran  0.005ns 3ns

.control
  run
  * >>>>> plot >>>>>>
  set xgridwidth  = 2
  set xbrushwidth = 3
  * "svgwidth", "svgheight",  "svgfont-size", "svgfont-width", "svguse-color", "svgstroke-width", "svggrid-width",
  set svg_intopts = ( 1024 256 16 0 1 2 0 )
  * "svgbackground", "svgfont-family", "svgfont"
  setcs svg_stropts = ( white Arial Arial )
  set hcopydevtype = svg
  set color1       = black
  set color2       = red
  set color3       = blue
  set color4       = green

  hardcopy fig/plot_and8c_t.svg
  + in1 out in8
  + title 'CMOS AND8c'
  + xlabel 't'
  + ylabel 'Voltage'
  + ylimit 0 1.5
  + ydelta 0.5

  * for MS Windows, using Edge
  if $oscompiled = 1 | $oscompiled = 8
    shell Start fig/plot_and8c_t.svg
  else
    if $oscompiled = 7
      * macOS (using Safari, no need to install X11)
      shell open -a safari fig/plot_and8c_t.svg &
    else
      * for CYGWIN, Linux, using feh and X11
      shell feh --magick-timeout 1 fig/plot_and8c_t.svg &
    end
  end
  * <<<<< plot <<<<<
.endc

* Measurement
* -----------------------------------------------------------------------------
.measure tran tr   trig V(out) val='VDD*0.1' rise=1 targ V(out) val='VDD*0.9' rise=1
.measure tran tf   trig V(out) val='VDD*0.9' fall=1 targ V(out) val='VDD*0.1' fall=1
.measure tran tpdr trig V(in1) val='VDD/2'   rise=1 targ V(out) val='VDD/2'   rise=1
.measure tran tpdf trig V(in8) val='VDD/2'   fall=1 targ V(out) val='VDD/2'   fall=1
.measure tran tpd  param='(tpdr+tpdf)/2'

* power dissipation of the AND8 gate
.inc ./and8_test_pow.inc

.end
